library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package FIR_package IS
    type Taps_array is array (natural range 0 to 10) of std_logic_vector(15 downto 0);
	 type MAC_array is array (natural range 0 to 10) of std_logic_vector(31 downto 0);
	 type Coeffs_array is array (natural range 0 to 10) of std_logic_vector(15 downto 0);
end package; 